//
// File: top_pkg.sv
//
// Generated from Mentor VIP Configurator (20210701)
// Generated using Mentor VIP Library ( 2021.3_2 : 09/26/2021:08:26 )
//
package top_pkg;
    import uvm_pkg::*;
    
    `include "uvm_macros.svh"
    
    import addr_map_pkg::*;
    
    import top_params_pkg::*;
    import mvc_pkg::*;
    import mgc_axi4lite_seq_pkg::*;
    import mgc_axi4_v1_0_pkg::*;
    
    `include "top_env_config.svh"
    `include "top_env.svh"
    `include "top_vseq_base.svh"
    `include "top_test_base.svh"
    `include "top_example_vseq.svh"
endpackage: top_pkg
