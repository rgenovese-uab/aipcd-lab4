//
// File: test_packages.svh
//
// Generated from Mentor VIP Configurator (20210701)
// Generated using Mentor VIP Library ( 2021.3_2 : 09/26/2021:08:26 )
//

import top_pkg::*;

// Add other packages here as required
